// iHCF Configuration File
// This is in a new custom format **NOT YAML**
// Be sure to double-check your config
// Credits - Techcable's Configuration API

// If the plugin should attempt to limit entities to reduce lag.
// currently what this does is allow only 25 entities in one chunk.
handleEntityLimiting = true

// If arrows shot from a bow with infinity should be removed
// when they land to reduce entity lag.
removeInfinityArrowsOnLand = true

// The maximum Beacon strength level
beaconStrengthLevelLimit = 1

// If boats should not be allowed to be placed on land.
disableBoatPlacementOnLand = true

enderpearlGlitching {
     // If this plugin should try and block Enderpearl glitching.
     enabled = true

     // If the enderpearl should be refunded if the player was detected.
     refund = true
}

// If enderchests should be disabled.
disableEnderchests = true

// If beds cannot be placed in the Nether.
preventPlacingBedsNether = true

// Timezone to use for events and stuff
serverTimeZone = EST

// The speed at which items in furnaces cook, set to 1.0 for default.
furnaceCookSpeedMultiplier = 6.0

// If you should be able to bottle exp by crafting a glass bottle.
bottledExp = true

// If you should be able to de-enchant books by right clicking enchant tables.
bookDeenchanting = true

// If death signs should spawn upon deaths.
deathSigns = true

// If death signs should thaw upon deaths.
deathLightning = true

// The current number of the map.
mapNumber = 1

// If the server is in a kit map mode.
kitMap = false

// If ally damage should be prevented or just warn the attacker.
preventAllyDamage = true

economy {
    // The amount of money a player starts off with.
    startingBalance = 250
}

spawners {
    // If players should not be able to break spawners in the Nether.
    preventBreakingNether = true

    // If players should not be able to place spawners in the Nether.
    preventPlacingNether = true
}

expMultiplier {
    // The multipliers to set for experience, set to 1.0 to normalise as vanilla.
    global = 2.0
    fishing = 2.0
    smelting = 2.0
    lootingPerLevel = 1.5
    luckPerLevel = 1.5
    fortunePerLevel = 1.5
}

scoreboard {
    sidebar {
        // The title of the sidebar, use {MAP_NUMBER} as a
        // placeholder with & as colour codes.
        title = "&a&lHCF &c[Map {MAP_NUMBER}]"

        // If this plugin utilises the sidebar.
        enabled = true

        // All scoreboard entries must be below 48 characters,
        // including color codes (-> &e15 characters <-).  Please
        // keep note of your maximum faction character limit.
        eotw {

        }
    }

    tablist {
        // Custom Tablist
        title = "&a&lHCF"

        // If this plugin utilizes the custom tablist.
        enabled = true
    }

    nametags {
        // If this plugin will utilise nametags.
        enabled = true
    }
}

combatlog {
    // If this plugin will protect from combat-logging.
    enabled = true

    // The ticks for when a combat logger NPC should despawn.
    despawnDelayTicks = 600
}

warzone {
    // The radius of the warzone.
    radiusOverworld = 800
    radiusNether = 800
}

factions {
    conquest {
        // How much points should a faction lose when a player dies in Conquest.
        pointLossPerDeath = 20

        // How much points should a faction need to win Conquest.
        requiredVictoryPoints = 300

        // If negative points are possible during conquest.
        allowNegativePoints = true
    }

    roads {
        // If players are allowed to claim next to roads
        allowClaimsBesides = true
    }

    // List of faction names that cannot be used.
    disallowedFactionNames = [
        "EOTW",
        "KOHI"
    ]

    home {
        // The time in seconds to teleport to faction home, -1 to disable, 0 for instant
        teleportDelay {
            NETHER = 30
            THE_END = -1
            NORMAL = 10
        }

        // The maximum height to set a faction home, use -1 to ignore this.
        maxHeight = -1

        // If faction homing in enemy territory should be allowed.
        allowTeleportingInEnemyTerritory = true
    }

    // Minimum amount of characters a faction name must be.
    nameMinCharacters = 3

    // Maximum amount of characters a faction name must be.
    nameMaxCharacters = 16

    // Maximum amount of members a faction can own.
    maxMembers = 25

    // Maximum amount of claims a faction can own.
    maxClaims = 8

    // Maximum amount of allies a faction can have.
    maxAllies = 1

    subclaim {
        // The minimum characters a player can name a subclaim.
        nameMinCharacters = 3

        // The maximum characters a player can name a subclaim.
        nameMaxCharacters = 16
    }

    dtr {
        regenFreeze {
            // The minutes for faction DTR regen freeze to
            // end not including any multipliers, etc.
            baseMinutes = 40

            // How much longer the DTR freeze should be for factions with
            // more members. Set to 0 to disable.
            minutesPerMember = 2
        }

        // The minimum DTR a faction can have.
        minimum = -50

        // The maximum DTR a faction will regenerate to.
        maximum = 6

        // Time in milliseconds between a DTR update.
        millisecondsBetweenUpdates = 45000

        // The DTR again when DTR updates.
        incrementBetweenUpdates = 0.1
    }

    relationColours {
        // The nametag and chat colours to show for faction relations.
        wilderness = "DARK_GREEN"
        warzone = "LIGHT_PURPLE"
        teammate = "GREEN"
        ally = "GOLD"
        enemy = "RED"
        road = "YELLOW"
        safezone = "AQUA"
    }
}

deathban {
    // The regular deathban duration.
    baseDurationMinutes = 60

    // The seconds before kicking after showing the user
    // the respawn screen from a deathban.
    respawnScreenSecondsBeforeKick = 15
}

end {
    // If the end should be opened.
    open = true

    // The location of the spawn point when leaving end by End Portal.
    exitLocation = "world,0.5,75,0.5,0,0"

    // If fire should be extinguished when leaving the end through an End Portal.
    extinguishFireOnExit = true

    // If strength should be removed when entering the end through an End Portal.
    removeStrengthOnEntrance = true
}

eotw {
    chatSymbolPrefix = " \u2605"
    chatSymbolSuffix = ""

    // List of UUIDs that capped last maps EOTW.
    lastMapCapperUuids = [
    ]
}

// The maximum levels an enchantment can be.
enchantmentLimits = [
    "PROTECTION_ENVIRONMENTAL = 3",
    "PROTECTION_FIRE = 3",
    "SILK_TOUCH = 1",
    "DURABILITY = 3",
    "PROTECTION_EXPLOSIONS = 3",
    "LOOT_BONUS_BLOCKS = 3",
    "PROTECTION_PROJECTILE = 3",
    "OXYGEN = 3",
    "WATER_WORKER = 1",
    "THORNS = 0",
    "DAMAGE_ALL = 3",
    "ARROW_KNOCKBACK = 1",
    "KNOCKBACK = 1",
    "FIRE_ASPECT = 1",
    "LOOT_BONUS_MOBS = 3",
    "LUCK = 3",
    "LURE = 3",
    "DEPTH_STRIDER = 0"
]

// The maximum levels a potion can be brewed to.
potionLimits = [
    "STRENGTH = 0",
    "INVISIBILITY = 0",
    "REGEN = 0",
    "WEAKNESS = 0",
    "INSTANT_DAMAGE = 0",
    "SLOWNESS = 1",
    "POISON = 1"
]

subclaimSigns {
    // Protects against members that are not on the sign opening.
    private = false

    // Protects against any non-officer opening.
    captain = true

    // Protects against any non-leader opening.
    leader = false

    // If subclaim protected objects should be protected from hopper
    // items too, disabling this may increase performance.
    hopperCheck = true
}